module lab2(a,e);

input [3:0] a;
output [6:0] e;

//0
assign e[6] =(~a[3]&~a[2]&~a[1]&a[0])|(~a[3]&a[2]&~a[1]&~a[0])|(a[3]&~a[2]&a[1]&a[0])|(a[3]&a[2]&~a[1]&a[0]);
//1
assign e[5] = (~a[3]&a[2]&~a[1]&a[0])|(a[2]&a[1]&~a[0])|(a[3]&a[2]&~a[0])|(a[3]&a[1]&a[0]);

//2
assign e[4]= (~a[3]&~a[2]&a[1]&~a[0])|(a[3]&a[2]&~a[0])|(a[3]&a[2]&a[1]);

//3
assign e[3]= (~a[3]&~a[2]&~a[1]&a[0])|(~a[3]&a[2]&~a[1]&~a[0])|(a[3]&~a[2]&a[1]&~a[0])|(a[2]&a[1]&a[0]);
//4
assign e[2]= (~a[2]&~a[1]&a[0])|(~a[3]&a[2]&~a[1])|(~a[3]&a[0]);
//5
assign e[1]= (a[3]&a[2]&~a[1]&a[0])|(~a[3]&~a[2]&a[0])|(~a[3]&~a[2]&a[1])|(~a[3]&a[1]&a[0]);

//6


// In minterm form, the function was originally f = ~a[3]~a[2]~a[1]~a[0] + ~a[3]~a[2]~a[1]~a[0] + ~a[3]a[2]a[1]a[0] + a[3]a[2]~a[1]~a[0]

// f = ~a[3]~a[2]~a[1]~a[0] + ~a[3]~a[2]~a[1]a[0] + ~a[3]a[2]a[1]a[0] + a[3]a[2]~a[1]~a[0]

// = ~a[3]~a[2]~a[1](~a[0] + a[0]) + ~a[3]a[2]a[1]a[0] + a[3]a[2]~a[1]~a[0]

// = ~a[3]~a[2]~a[1](1) + ~a[3]a[2]a[1]a[0] + a[3]a[2]~a[1]~a[0]


assign e[0]= (~a[3]&a[2]&a[1]&a[0])|(a[3]&a[2]&~a[1]&~a[0])|(~a[3]&~a[2]&~a[1]);

endmodule