//module remove2complement(a, f);
//
//input [3:0] a;
//
//output[3:0] f;
//wire cout;
//
//wire [3:0] int;
//
//assign int[0] = ~a[0];
//assign int[1] = ~a[1];
//assign int[2] = ~a[2];
//assign int[3] = ~a[3];
//
//ripplecarry(int, 0001, 0, f, cout);
//
////assign g = cout + ~op;
//
//endmodule
